module TopModule(input sw, output led);
	assign led = sw;
endmodule